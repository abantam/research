module sp_build_bv #(
	parameter num_of_rules = 1000
)(
	input  clk,rst,
	input  [num_of_rules:0] rules,
	output [31:0] match_bv
);

initial begin
	
end

endmodule
