// unsaved.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module unsaved (
		input  wire         clk_clk,                           //                     clk.clk
		output wire         clk_0_clk_clk,                     //               clk_0_clk.clk
		output wire         clk_0_clk_reset_reset_n,           //         clk_0_clk_reset.reset_n
		input  wire         onchip_memory2_0_clk1_clk,         //   onchip_memory2_0_clk1.clk
		input  wire         onchip_memory2_0_reset1_reset,     // onchip_memory2_0_reset1.reset
		input  wire         onchip_memory2_0_reset1_reset_req, //                        .reset_req
		input  wire [7:0]   onchip_memory2_0_s1_address,       //     onchip_memory2_0_s1.address
		input  wire         onchip_memory2_0_s1_clken,         //                        .clken
		input  wire         onchip_memory2_0_s1_chipselect,    //                        .chipselect
		input  wire         onchip_memory2_0_s1_write,         //                        .write
		output wire [127:0] onchip_memory2_0_s1_readdata,      //                        .readdata
		input  wire [127:0] onchip_memory2_0_s1_writedata,     //                        .writedata
		input  wire [15:0]  onchip_memory2_0_s1_byteenable,    //                        .byteenable
		input  wire         reset_reset_n                      //                   reset.reset_n
	);

	unsaved_onchip_memory2_0 onchip_memory2_0 (
		.clk        (onchip_memory2_0_clk1_clk),         //   clk1.clk
		.address    (onchip_memory2_0_s1_address),       //     s1.address
		.clken      (onchip_memory2_0_s1_clken),         //       .clken
		.chipselect (onchip_memory2_0_s1_chipselect),    //       .chipselect
		.write      (onchip_memory2_0_s1_write),         //       .write
		.readdata   (onchip_memory2_0_s1_readdata),      //       .readdata
		.writedata  (onchip_memory2_0_s1_writedata),     //       .writedata
		.byteenable (onchip_memory2_0_s1_byteenable),    //       .byteenable
		.reset      (onchip_memory2_0_reset1_reset),     // reset1.reset
		.reset_req  (onchip_memory2_0_reset1_reset_req)  //       .reset_req
	);

	assign clk_0_clk_clk = clk_clk;

	assign clk_0_clk_reset_reset_n = reset_reset_n;

endmodule
