module FSBV(
	input  clk,rst,
	input  [103:0] pkt_header,
	output [31:0] matching_bv
);

parameter num_of_rules = 1000;

endmodule