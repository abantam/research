module sp_build_bv #(
	parameter num_of_rules = 10
)(
	input  clk,rst,
	input  [num_of_rules-1:0] rules,
	output [31:0] match_bv
);

initial begin
	
end

endmodule
