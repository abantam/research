module gen_bit_vector(
	
);

endmodule