module openflow13(
	input [10:0] packet,
	output [10:0] bit_vector
);

endmodule